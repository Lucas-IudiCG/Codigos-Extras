<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-3.85,35.1565,83.35,-61.5101</PageViewport>
<gate>
<ID>2</ID>
<type>AI_XOR2</type>
<position>16.5,-26</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>1 </input>
<output>
<ID>OUT</ID>3 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4</ID>
<type>AI_XOR2</type>
<position>28.5,-26</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>1 </input>
<output>
<ID>OUT</ID>4 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6</ID>
<type>AI_XOR2</type>
<position>40.5,-26</position>
<input>
<ID>IN_0</ID>14 </input>
<input>
<ID>IN_1</ID>1 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8</ID>
<type>AI_XOR2</type>
<position>53,-26</position>
<input>
<ID>IN_0</ID>20 </input>
<input>
<ID>IN_1</ID>1 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_TOGGLE</type>
<position>71.5,-32</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_TOGGLE</type>
<position>17.5,-8.5</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_TOGGLE</type>
<position>22.5,-8.5</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_FULLADDER_1BIT</type>
<position>17.5,-32</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_B_0</ID>3 </input>
<output>
<ID>OUT_0</ID>16 </output>
<input>
<ID>carry_in</ID>5 </input>
<output>
<ID>carry_out</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_FULLADDER_1BIT</type>
<position>29.5,-32</position>
<input>
<ID>IN_0</ID>13 </input>
<input>
<ID>IN_B_0</ID>4 </input>
<output>
<ID>OUT_0</ID>17 </output>
<input>
<ID>carry_in</ID>8 </input>
<output>
<ID>carry_out</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>20</ID>
<type>GA_LED</type>
<position>8,-38</position>
<input>
<ID>N_in3</ID>11 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>22</ID>
<type>GA_LED</type>
<position>17.5,-38</position>
<input>
<ID>N_in3</ID>16 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>GA_LED</type>
<position>29.5,-38</position>
<input>
<ID>N_in3</ID>17 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>26</ID>
<type>GA_LED</type>
<position>41.5,-38</position>
<input>
<ID>N_in3</ID>18 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>28</ID>
<type>GA_LED</type>
<position>54,-38</position>
<input>
<ID>N_in3</ID>19 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>30</ID>
<type>AA_FULLADDER_1BIT</type>
<position>41.5,-32</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_B_0</ID>7 </input>
<output>
<ID>OUT_0</ID>18 </output>
<input>
<ID>carry_in</ID>10 </input>
<output>
<ID>carry_out</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>32</ID>
<type>AA_FULLADDER_1BIT</type>
<position>54,-32</position>
<input>
<ID>IN_0</ID>21 </input>
<input>
<ID>IN_B_0</ID>9 </input>
<output>
<ID>OUT_0</ID>19 </output>
<input>
<ID>carry_in</ID>1 </input>
<output>
<ID>carry_out</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>34</ID>
<type>AA_TOGGLE</type>
<position>29.5,-8.5</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>36</ID>
<type>AA_TOGGLE</type>
<position>34,-8.5</position>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>38</ID>
<type>AA_TOGGLE</type>
<position>41.5,-8.5</position>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>40</ID>
<type>AA_TOGGLE</type>
<position>46.5,-8.5</position>
<output>
<ID>OUT_0</ID>15 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>42</ID>
<type>AA_TOGGLE</type>
<position>59,-8.5</position>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_TOGGLE</type>
<position>54.5,-8.5</position>
<output>
<ID>OUT_0</ID>20 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>46</ID>
<type>AA_LABEL</type>
<position>17,-5</position>
<gparam>LABEL_TEXT B3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>48</ID>
<type>AA_LABEL</type>
<position>23,-5.5</position>
<gparam>LABEL_TEXT A3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>50</ID>
<type>AA_LABEL</type>
<position>29,-5</position>
<gparam>LABEL_TEXT B2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>52</ID>
<type>AA_LABEL</type>
<position>34,-5</position>
<gparam>LABEL_TEXT A2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>54</ID>
<type>AA_LABEL</type>
<position>41.5,-5</position>
<gparam>LABEL_TEXT B1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>56</ID>
<type>AA_LABEL</type>
<position>47,-5</position>
<gparam>LABEL_TEXT A1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>58</ID>
<type>AA_LABEL</type>
<position>55,-4.5</position>
<gparam>LABEL_TEXT B0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>60</ID>
<type>AA_LABEL</type>
<position>59,-5</position>
<gparam>LABEL_TEXT A0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>62</ID>
<type>AA_LABEL</type>
<position>71.5,-28</position>
<gparam>LABEL_TEXT Te</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>64</ID>
<type>AA_LABEL</type>
<position>8,-42</position>
<gparam>LABEL_TEXT S4</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>66</ID>
<type>AA_LABEL</type>
<position>17.5,-42</position>
<gparam>LABEL_TEXT S3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>68</ID>
<type>AA_LABEL</type>
<position>29.5,-41.5</position>
<gparam>LABEL_TEXT S2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>70</ID>
<type>AA_LABEL</type>
<position>41,-41.5</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>72</ID>
<type>AA_LABEL</type>
<position>54,-41.5</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15.5,-23,15.5,-14</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>-14 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15.5,-14,65,-14</points>
<intersection>15.5 0</intersection>
<intersection>27.5 4</intersection>
<intersection>39.5 5</intersection>
<intersection>52 6</intersection>
<intersection>65 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>65,-32,65,-14</points>
<intersection>-32 3</intersection>
<intersection>-14 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>58,-32,69.5,-32</points>
<connection>
<GID>32</GID>
<name>carry_in</name></connection>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>65 2</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>27.5,-23,27.5,-14</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<intersection>-14 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>39.5,-23,39.5,-14</points>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<intersection>-14 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>52,-23,52,-14</points>
<connection>
<GID>8</GID>
<name>IN_1</name></connection>
<intersection>-14 1</intersection></vsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17.5,-23,17.5,-10.5</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<intersection>-23 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>17.5,-23,17.5,-23</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>17.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16.5,-29,16.5,-29</points>
<connection>
<GID>2</GID>
<name>OUT</name></connection>
<connection>
<GID>16</GID>
<name>IN_B_0</name></connection></vsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,-29,28.5,-29</points>
<connection>
<GID>18</GID>
<name>IN_B_0</name></connection>
<connection>
<GID>4</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>21.5,-32,25.5,-32</points>
<connection>
<GID>16</GID>
<name>carry_in</name></connection>
<connection>
<GID>18</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18.5,-29,18.5,-27.5</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>-27.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>22.5,-27.5,22.5,-10.5</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>-27.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>18.5,-27.5,22.5,-27.5</points>
<intersection>18.5 0</intersection>
<intersection>22.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,-29,40.5,-29</points>
<connection>
<GID>6</GID>
<name>OUT</name></connection>
<connection>
<GID>30</GID>
<name>IN_B_0</name></connection></vsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>33.5,-32,37.5,-32</points>
<connection>
<GID>18</GID>
<name>carry_in</name></connection>
<connection>
<GID>30</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53,-29,53,-29</points>
<connection>
<GID>8</GID>
<name>OUT</name></connection>
<connection>
<GID>32</GID>
<name>IN_B_0</name></connection></vsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-32,50,-32</points>
<connection>
<GID>30</GID>
<name>carry_in</name></connection>
<connection>
<GID>32</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8,-37,8,-32</points>
<connection>
<GID>20</GID>
<name>N_in3</name></connection>
<intersection>-32 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>8,-32,13.5,-32</points>
<connection>
<GID>16</GID>
<name>carry_out</name></connection>
<intersection>8 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29.5,-23,29.5,-10.5</points>
<connection>
<GID>34</GID>
<name>OUT_0</name></connection>
<intersection>-23 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>29.5,-23,29.5,-23</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>29.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-27.5,34,-10.5</points>
<connection>
<GID>36</GID>
<name>OUT_0</name></connection>
<intersection>-27.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>30.5,-29,30.5,-27.5</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>-27.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>30.5,-27.5,34,-27.5</points>
<intersection>30.5 1</intersection>
<intersection>34 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41.5,-23,41.5,-10.5</points>
<connection>
<GID>38</GID>
<name>OUT_0</name></connection>
<intersection>-23 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>41.5,-23,41.5,-23</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>41.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42.5,-29,42.5,-28</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<intersection>-28 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>46.5,-28,46.5,-10.5</points>
<connection>
<GID>40</GID>
<name>OUT_0</name></connection>
<intersection>-28 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>42.5,-28,46.5,-28</points>
<intersection>42.5 0</intersection>
<intersection>46.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17.5,-37,17.5,-35</points>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection>
<connection>
<GID>22</GID>
<name>N_in3</name></connection></vsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29.5,-37,29.5,-35</points>
<connection>
<GID>24</GID>
<name>N_in3</name></connection>
<connection>
<GID>18</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41.5,-37,41.5,-35</points>
<connection>
<GID>26</GID>
<name>N_in3</name></connection>
<connection>
<GID>30</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,-37,54,-35</points>
<connection>
<GID>32</GID>
<name>OUT_0</name></connection>
<connection>
<GID>28</GID>
<name>N_in3</name></connection></vsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,-23,54.5,-10.5</points>
<connection>
<GID>44</GID>
<name>OUT_0</name></connection>
<intersection>-23 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>54,-23,54.5,-23</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>54.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55,-29,55,-27.5</points>
<connection>
<GID>32</GID>
<name>IN_0</name></connection>
<intersection>-27.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>59,-27.5,59,-10.5</points>
<connection>
<GID>42</GID>
<name>OUT_0</name></connection>
<intersection>-27.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>55,-27.5,59,-27.5</points>
<intersection>55 0</intersection>
<intersection>59 1</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,65.4,-72.5</PageViewport></page 1>
<page 2>
<PageViewport>0,0,65.4,-72.5</PageViewport></page 2>
<page 3>
<PageViewport>0,0,65.4,-72.5</PageViewport></page 3>
<page 4>
<PageViewport>0,0,65.4,-72.5</PageViewport></page 4>
<page 5>
<PageViewport>0,0,65.4,-72.5</PageViewport></page 5>
<page 6>
<PageViewport>0,0,65.4,-72.5</PageViewport></page 6>
<page 7>
<PageViewport>0,0,65.4,-72.5</PageViewport></page 7>
<page 8>
<PageViewport>0,0,65.4,-72.5</PageViewport></page 8>
<page 9>
<PageViewport>0,0,65.4,-72.5</PageViewport></page 9></circuit>