<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-42.5789,75.0501,194.488,-47.2166</PageViewport>
<gate>
<ID>2</ID>
<type>AA_AND2</type>
<position>21,-7.5</position>
<input>
<ID>IN_0</ID>14 </input>
<input>
<ID>IN_1</ID>16 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4</ID>
<type>BE_NOR2</type>
<position>23,-52</position>
<input>
<ID>IN_0</ID>14 </input>
<input>
<ID>IN_1</ID>16 </input>
<output>
<ID>OUT</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6</ID>
<type>BA_NAND2</type>
<position>22,-36</position>
<input>
<ID>IN_0</ID>14 </input>
<input>
<ID>IN_1</ID>16 </input>
<output>
<ID>OUT</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8</ID>
<type>AE_OR2</type>
<position>22,-22</position>
<input>
<ID>IN_0</ID>14 </input>
<input>
<ID>IN_1</ID>16 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>10</ID>
<type>GA_LED</type>
<position>53,-7.5</position>
<input>
<ID>N_in0</ID>7 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>GA_LED</type>
<position>53,-16</position>
<input>
<ID>N_in0</ID>5 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>14</ID>
<type>BE_NOR2</type>
<position>22.5,-16</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>16</ID>
<type>BA_NAND2</type>
<position>22,-29</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>4 </input>
<output>
<ID>OUT</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>18</ID>
<type>BI_NANDX2</type>
<position>22.5,-43.5</position>
<input>
<ID>IN_0</ID>14 </input>
<input>
<ID>IN_1</ID>16 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>20</ID>
<type>BM_NORX2</type>
<position>22.5,-59</position>
<input>
<ID>IN_0</ID>14 </input>
<input>
<ID>IN_1</ID>16 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>22</ID>
<type>AE_SMALL_INVERTER</type>
<position>17.5,-15</position>
<input>
<ID>IN_0</ID>14 </input>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>24</ID>
<type>AE_SMALL_INVERTER</type>
<position>17.5,-17</position>
<input>
<ID>IN_0</ID>16 </input>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>26</ID>
<type>AE_SMALL_INVERTER</type>
<position>17,-28</position>
<input>
<ID>IN_0</ID>14 </input>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>28</ID>
<type>AE_SMALL_INVERTER</type>
<position>17,-30</position>
<input>
<ID>IN_0</ID>16 </input>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>30</ID>
<type>GA_LED</type>
<position>53.5,-22</position>
<input>
<ID>N_in0</ID>8 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>32</ID>
<type>GA_LED</type>
<position>53.5,-29</position>
<input>
<ID>N_in0</ID>13 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>GA_LED</type>
<position>54,-36</position>
<input>
<ID>N_in0</ID>12 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>36</ID>
<type>GA_LED</type>
<position>54,-43.5</position>
<input>
<ID>N_in0</ID>11 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>38</ID>
<type>GA_LED</type>
<position>54,-51.5</position>
<input>
<ID>N_in0</ID>10 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>40</ID>
<type>GA_LED</type>
<position>54,-59</position>
<input>
<ID>N_in0</ID>9 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>42</ID>
<type>AA_TOGGLE</type>
<position>-28,-20</position>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_TOGGLE</type>
<position>-28.5,-35</position>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>46</ID>
<type>AA_LABEL</type>
<position>-27.5,-15</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>48</ID>
<type>AA_LABEL</type>
<position>-28.5,-30.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>50</ID>
<type>AA_LABEL</type>
<position>53,-4.5</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>52</ID>
<type>AA_LABEL</type>
<position>53,-13</position>
<gparam>LABEL_TEXT 2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>54</ID>
<type>AA_LABEL</type>
<position>53.5,-19.5</position>
<gparam>LABEL_TEXT 3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>56</ID>
<type>AA_LABEL</type>
<position>53,-25.5</position>
<gparam>LABEL_TEXT 4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>58</ID>
<type>AA_LABEL</type>
<position>53.5,-33.5</position>
<gparam>LABEL_TEXT 5</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>60</ID>
<type>AA_LABEL</type>
<position>53.5,-41</position>
<gparam>LABEL_TEXT 6</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>62</ID>
<type>AA_LABEL</type>
<position>54,-48.5</position>
<gparam>LABEL_TEXT 7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>64</ID>
<type>AA_LABEL</type>
<position>54,-56</position>
<gparam>LABEL_TEXT 8</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>66</ID>
<type>AA_LABEL</type>
<position>12.5,33</position>
<gparam>LABEL_TEXT Exercicio 3.1.2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19.5,-15,19.5,-15</points>
<connection>
<GID>22</GID>
<name>OUT_0</name></connection>
<connection>
<GID>14</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19.5,-17,19.5,-17</points>
<connection>
<GID>14</GID>
<name>IN_1</name></connection>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19,-28,19,-28</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<connection>
<GID>16</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19,-30,19,-30</points>
<connection>
<GID>16</GID>
<name>IN_1</name></connection>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25.5,-16,52,-16</points>
<connection>
<GID>14</GID>
<name>OUT</name></connection>
<connection>
<GID>12</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24,-7.5,52,-7.5</points>
<connection>
<GID>2</GID>
<name>OUT</name></connection>
<connection>
<GID>10</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25,-22,52.5,-22</points>
<connection>
<GID>30</GID>
<name>N_in0</name></connection>
<connection>
<GID>8</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25.5,-59,53,-59</points>
<connection>
<GID>20</GID>
<name>OUT</name></connection>
<connection>
<GID>40</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26,-52,53,-52</points>
<connection>
<GID>4</GID>
<name>OUT</name></connection>
<intersection>53 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>53,-52,53,-51.5</points>
<connection>
<GID>38</GID>
<name>N_in0</name></connection>
<intersection>-52 1</intersection></vsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25.5,-43.5,53,-43.5</points>
<connection>
<GID>18</GID>
<name>OUT</name></connection>
<connection>
<GID>36</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25,-36,53,-36</points>
<connection>
<GID>34</GID>
<name>N_in0</name></connection>
<connection>
<GID>6</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25,-29,52.5,-29</points>
<connection>
<GID>16</GID>
<name>OUT</name></connection>
<connection>
<GID>32</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>4,-58,4,-6.5</points>
<intersection>-58 11</intersection>
<intersection>-51 8</intersection>
<intersection>-42.5 12</intersection>
<intersection>-35 6</intersection>
<intersection>-28 10</intersection>
<intersection>-21 14</intersection>
<intersection>-20 2</intersection>
<intersection>-15 4</intersection>
<intersection>-6.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>4,-6.5,18,-6.5</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>4 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-26,-20,4,-20</points>
<connection>
<GID>42</GID>
<name>OUT_0</name></connection>
<intersection>4 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>4,-15,15.5,-15</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>4 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>4,-35,19,-35</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>4 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>4,-51,20,-51</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>4 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>4,-28,15,-28</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>4 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>4,-58,19.5,-58</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>4 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>4,-42.5,19.5,-42.5</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>4 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>4,-21,19,-21</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>4 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4,-60,-4,-8.5</points>
<intersection>-60 9</intersection>
<intersection>-53 11</intersection>
<intersection>-44.5 7</intersection>
<intersection>-37 10</intersection>
<intersection>-35 2</intersection>
<intersection>-30 4</intersection>
<intersection>-23 13</intersection>
<intersection>-17 5</intersection>
<intersection>-8.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4,-8.5,18,-8.5</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>-4 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-26.5,-35,-4,-35</points>
<connection>
<GID>44</GID>
<name>OUT_0</name></connection>
<intersection>-4 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-4,-30,15,-30</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<intersection>-4 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-4,-17,15.5,-17</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>-4 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-4,-44.5,19.5,-44.5</points>
<connection>
<GID>18</GID>
<name>IN_1</name></connection>
<intersection>-4 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-4,-60,19.5,-60</points>
<connection>
<GID>20</GID>
<name>IN_1</name></connection>
<intersection>-4 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-4,-37,19,-37</points>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<intersection>-4 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-4,-53,20,-53</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<intersection>-4 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-4,-23,19,-23</points>
<connection>
<GID>8</GID>
<name>IN_1</name></connection>
<intersection>-4 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,177.8,-91.7</PageViewport></page 1>
<page 2>
<PageViewport>0,0,177.8,-91.7</PageViewport></page 2>
<page 3>
<PageViewport>0,0,177.8,-91.7</PageViewport></page 3>
<page 4>
<PageViewport>0,0,177.8,-91.7</PageViewport></page 4>
<page 5>
<PageViewport>0,0,177.8,-91.7</PageViewport></page 5>
<page 6>
<PageViewport>0,0,177.8,-91.7</PageViewport></page 6>
<page 7>
<PageViewport>0,0,177.8,-91.7</PageViewport></page 7>
<page 8>
<PageViewport>0,0,177.8,-91.7</PageViewport></page 8>
<page 9>
<PageViewport>0,0,177.8,-91.7</PageViewport></page 9></circuit>