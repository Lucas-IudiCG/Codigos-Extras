<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-16.4,11.7333,66.8,-82.1333</PageViewport>
<gate>
<ID>2</ID>
<type>AA_TOGGLE</type>
<position>-8,-2.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>0,-6</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>-7.5,-21</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_TOGGLE</type>
<position>-7.5,-27</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_AND2</type>
<position>16,-3.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_AND2</type>
<position>14,-17.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>7 </input>
<output>
<ID>OUT</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>14</ID>
<type>AE_OR2</type>
<position>28,-9</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>16</ID>
<type>AE_OR2</type>
<position>2.5,-23.5</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_LABEL</type>
<position>-7,0.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>AA_LABEL</type>
<position>1,-3.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>22</ID>
<type>AA_LABEL</type>
<position>-7.5,-19</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>AA_LABEL</type>
<position>-7.5,-23.5</position>
<gparam>LABEL_TEXT D</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>26</ID>
<type>GA_LED</type>
<position>32,-9</position>
<input>
<ID>N_in0</ID>8 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-2.5,-16.5,-2.5,-2.5</points>
<intersection>-16.5 4</intersection>
<intersection>-2.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-6,-2.5,13,-2.5</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>-2.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-2.5,-16.5,11,-16.5</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>-2.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5.5,-6,5.5,-4.5</points>
<intersection>-6 2</intersection>
<intersection>-4.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>5.5,-4.5,13,-4.5</points>
<connection>
<GID>10</GID>
<name>IN_1</name></connection>
<intersection>5.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>2,-6,5.5,-6</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>5.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21.5,-17.5,21.5,-10</points>
<intersection>-17.5 2</intersection>
<intersection>-10 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21.5,-10,25,-10</points>
<connection>
<GID>14</GID>
<name>IN_1</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17,-17.5,21.5,-17.5</points>
<connection>
<GID>12</GID>
<name>OUT</name></connection>
<intersection>21.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22,-8,22,-3.5</points>
<intersection>-8 1</intersection>
<intersection>-3.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22,-8,25,-8</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>22 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>19,-3.5,22,-3.5</points>
<connection>
<GID>10</GID>
<name>OUT</name></connection>
<intersection>22 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-5.5,-21,-2.5,-21</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>-2.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-2.5,-22.5,-2.5,-21</points>
<intersection>-22.5 4</intersection>
<intersection>-21 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-2.5,-22.5,-0.5,-22.5</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>-2.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3,-27,-3,-24.5</points>
<intersection>-27 2</intersection>
<intersection>-24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-3,-24.5,-0.5,-24.5</points>
<connection>
<GID>16</GID>
<name>IN_1</name></connection>
<intersection>-3 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-5.5,-27,-3,-27</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>-3 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8,-23.5,8,-18.5</points>
<intersection>-23.5 2</intersection>
<intersection>-18.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>8,-18.5,11,-18.5</points>
<connection>
<GID>12</GID>
<name>IN_1</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>5.5,-23.5,8,-23.5</points>
<connection>
<GID>16</GID>
<name>OUT</name></connection>
<intersection>8 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,-9,31,-9</points>
<connection>
<GID>14</GID>
<name>OUT</name></connection>
<connection>
<GID>26</GID>
<name>N_in0</name></connection></vsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,62.4,-70.4</PageViewport></page 1>
<page 2>
<PageViewport>0,0,62.4,-70.4</PageViewport></page 2>
<page 3>
<PageViewport>0,0,62.4,-70.4</PageViewport></page 3>
<page 4>
<PageViewport>0,0,62.4,-70.4</PageViewport></page 4>
<page 5>
<PageViewport>0,0,62.4,-70.4</PageViewport></page 5>
<page 6>
<PageViewport>0,0,62.4,-70.4</PageViewport></page 6>
<page 7>
<PageViewport>0,0,62.4,-70.4</PageViewport></page 7>
<page 8>
<PageViewport>0,0,62.4,-70.4</PageViewport></page 8>
<page 9>
<PageViewport>0,0,62.4,-70.4</PageViewport></page 9></circuit>