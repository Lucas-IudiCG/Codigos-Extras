<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-3.18452e-006,0,93.6,-90.8</PageViewport>
<gate>
<ID>2</ID>
<type>AA_TOGGLE</type>
<position>8,-22.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>4</ID>
<type>BB_CLOCK</type>
<position>8,-27.5</position>
<output>
<ID>CLK</ID>2 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>8,-33.5</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_TOGGLE</type>
<position>8,-36</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_TOGGLE</type>
<position>8,-40.5</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_TOGGLE</type>
<position>8,-43</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>14</ID>
<type>DE_TO</type>
<position>18,-22.5</position>
<input>
<ID>IN_0</ID>1 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D</lparam></gate>
<gate>
<ID>16</ID>
<type>DE_TO</type>
<position>17.5,-27.5</position>
<input>
<ID>IN_0</ID>2 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CLK</lparam></gate>
<gate>
<ID>18</ID>
<type>DE_TO</type>
<position>18,-33.5</position>
<input>
<ID>IN_0</ID>3 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID J</lparam></gate>
<gate>
<ID>20</ID>
<type>DE_TO</type>
<position>18,-36</position>
<input>
<ID>IN_0</ID>4 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID K</lparam></gate>
<gate>
<ID>22</ID>
<type>DE_TO</type>
<position>17.5,-40.5</position>
<input>
<ID>IN_0</ID>5 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PR</lparam></gate>
<gate>
<ID>24</ID>
<type>DE_TO</type>
<position>17.5,-43</position>
<input>
<ID>IN_0</ID>6 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CLR</lparam></gate>
<gate>
<ID>26</ID>
<type>AE_DFF_LOW</type>
<position>61.5,-24.5</position>
<input>
<ID>IN_0</ID>13 </input>
<output>
<ID>OUTINV_0</ID>18 </output>
<output>
<ID>OUT_0</ID>17 </output>
<input>
<ID>clear</ID>11 </input>
<input>
<ID>clock</ID>14 </input>
<input>
<ID>set</ID>12 </input>
<gparam>angle 0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>30</ID>
<type>DA_FROM</type>
<position>61.5,-15.5</position>
<input>
<ID>IN_0</ID>12 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PR</lparam></gate>
<gate>
<ID>32</ID>
<type>DA_FROM</type>
<position>61.5,-32</position>
<input>
<ID>IN_0</ID>11 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID CLR</lparam></gate>
<gate>
<ID>34</ID>
<type>DA_FROM</type>
<position>61.5,-42.5</position>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PR</lparam></gate>
<gate>
<ID>36</ID>
<type>DA_FROM</type>
<position>61.5,-59</position>
<input>
<ID>IN_0</ID>23 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID CLR</lparam></gate>
<gate>
<ID>39</ID>
<type>DA_FROM</type>
<position>52,-22.5</position>
<input>
<ID>IN_0</ID>13 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D</lparam></gate>
<gate>
<ID>41</ID>
<type>DA_FROM</type>
<position>52,-25.5</position>
<input>
<ID>IN_0</ID>14 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CLK</lparam></gate>
<gate>
<ID>43</ID>
<type>DA_FROM</type>
<position>51.5,-45.5</position>
<input>
<ID>IN_0</ID>26 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID J</lparam></gate>
<gate>
<ID>45</ID>
<type>DA_FROM</type>
<position>51.5,-50</position>
<input>
<ID>IN_0</ID>25 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CLK</lparam></gate>
<gate>
<ID>47</ID>
<type>DE_TO</type>
<position>72.5,-22.5</position>
<input>
<ID>IN_0</ID>17 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID QD</lparam></gate>
<gate>
<ID>49</ID>
<type>DE_TO</type>
<position>72.5,-25.5</position>
<input>
<ID>IN_0</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID QD-</lparam></gate>
<gate>
<ID>51</ID>
<type>DE_TO</type>
<position>71.5,-48</position>
<input>
<ID>IN_0</ID>21 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID QJK</lparam></gate>
<gate>
<ID>53</ID>
<type>DE_TO</type>
<position>72,-52</position>
<input>
<ID>IN_0</ID>22 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID QJK-</lparam></gate>
<gate>
<ID>55</ID>
<type>DA_FROM</type>
<position>51.5,-54.5</position>
<input>
<ID>IN_0</ID>24 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID K</lparam></gate>
<gate>
<ID>57</ID>
<type>BE_JKFF_LOW</type>
<position>61.5,-50</position>
<input>
<ID>J</ID>26 </input>
<input>
<ID>K</ID>24 </input>
<output>
<ID>Q</ID>21 </output>
<input>
<ID>clear</ID>23 </input>
<input>
<ID>clock</ID>25 </input>
<output>
<ID>nQ</ID>22 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>10,-22.5,16,-22.5</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<connection>
<GID>14</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12,-27.5,15.5,-27.5</points>
<connection>
<GID>4</GID>
<name>CLK</name></connection>
<connection>
<GID>16</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>10,-33.5,16,-33.5</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<connection>
<GID>18</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>10,-36,16,-36</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<connection>
<GID>20</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>10,-40.5,15.5,-40.5</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<connection>
<GID>22</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>10,-43,15.5,-43</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<connection>
<GID>24</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61.5,-30,61.5,-28.5</points>
<connection>
<GID>26</GID>
<name>clear</name></connection>
<connection>
<GID>32</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61.5,-20.5,61.5,-17.5</points>
<connection>
<GID>26</GID>
<name>set</name></connection>
<connection>
<GID>30</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54,-22.5,58.5,-22.5</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<connection>
<GID>39</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54,-25.5,58.5,-25.5</points>
<connection>
<GID>26</GID>
<name>clock</name></connection>
<connection>
<GID>41</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>64.5,-22.5,70.5,-22.5</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<connection>
<GID>47</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>64.5,-25.5,70.5,-25.5</points>
<connection>
<GID>26</GID>
<name>OUTINV_0</name></connection>
<connection>
<GID>49</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>64.5,-48,69.5,-48</points>
<connection>
<GID>57</GID>
<name>Q</name></connection>
<connection>
<GID>51</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>64.5,-52,70,-52</points>
<connection>
<GID>57</GID>
<name>nQ</name></connection>
<connection>
<GID>53</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61.5,-57,61.5,-54</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<connection>
<GID>57</GID>
<name>clear</name></connection></vsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-54.5,56,-52</points>
<intersection>-54.5 2</intersection>
<intersection>-52 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56,-52,58.5,-52</points>
<connection>
<GID>57</GID>
<name>K</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>53.5,-54.5,56,-54.5</points>
<connection>
<GID>55</GID>
<name>IN_0</name></connection>
<intersection>56 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53.5,-50,58.5,-50</points>
<connection>
<GID>57</GID>
<name>clock</name></connection>
<connection>
<GID>45</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-48,56,-45.5</points>
<intersection>-48 1</intersection>
<intersection>-45.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56,-48,58.5,-48</points>
<connection>
<GID>57</GID>
<name>J</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>53.5,-45.5,56,-45.5</points>
<connection>
<GID>43</GID>
<name>IN_0</name></connection>
<intersection>56 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>20.475,-19.8625,73.125,-70.9375</PageViewport>
<gate>
<ID>3</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>68,-32</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>34 </input>
<input>
<ID>IN_2</ID>38 </input>
<input>
<ID>IN_3</ID>41 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 14</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>7</ID>
<type>GA_LED</type>
<position>25,-26</position>
<input>
<ID>N_in2</ID>41 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>11</ID>
<type>GA_LED</type>
<position>35.5,-26</position>
<input>
<ID>N_in2</ID>38 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>15</ID>
<type>GA_LED</type>
<position>46,-26.5</position>
<input>
<ID>N_in2</ID>34 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>19</ID>
<type>GA_LED</type>
<position>55.5,-26</position>
<input>
<ID>N_in2</ID>15 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>27</ID>
<type>AA_TOGGLE</type>
<position>9.5,-56</position>
<output>
<ID>OUT_0</ID>20 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>29</ID>
<type>AA_TOGGLE</type>
<position>9,-49.5</position>
<output>
<ID>OUT_0</ID>19 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>33</ID>
<type>AE_DFF_LOW</type>
<position>21.5,-42.5</position>
<input>
<ID>IN_0</ID>42 </input>
<output>
<ID>OUT_0</ID>41 </output>
<input>
<ID>clear</ID>20 </input>
<input>
<ID>clock</ID>19 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>37</ID>
<type>AE_DFF_LOW</type>
<position>31,-42.5</position>
<input>
<ID>IN_0</ID>41 </input>
<output>
<ID>OUT_0</ID>38 </output>
<input>
<ID>clear</ID>20 </input>
<input>
<ID>clock</ID>19 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>40</ID>
<type>AE_DFF_LOW</type>
<position>43,-42.5</position>
<input>
<ID>IN_0</ID>38 </input>
<output>
<ID>OUT_0</ID>34 </output>
<input>
<ID>clear</ID>20 </input>
<input>
<ID>clock</ID>19 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>44</ID>
<type>AE_DFF_LOW</type>
<position>51,-42.5</position>
<input>
<ID>IN_0</ID>34 </input>
<output>
<ID>OUT_0</ID>15 </output>
<input>
<ID>clear</ID>20 </input>
<input>
<ID>clock</ID>19 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>71</ID>
<type>AA_TOGGLE</type>
<position>9.5,-40.5</position>
<output>
<ID>OUT_0</ID>42 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>73</ID>
<type>AA_LABEL</type>
<position>8.5,-37</position>
<gparam>LABEL_TEXT Serial</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>75</ID>
<type>AA_LABEL</type>
<position>8.5,-53</position>
<gparam>LABEL_TEXT CLR</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>77</ID>
<type>AA_LABEL</type>
<position>8.5,-46</position>
<gparam>LABEL_TEXT CLK</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>79</ID>
<type>AA_LABEL</type>
<position>25,-23.5</position>
<gparam>LABEL_TEXT Q3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>81</ID>
<type>AA_LABEL</type>
<position>35,-23.5</position>
<gparam>LABEL_TEXT Q2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>83</ID>
<type>AA_LABEL</type>
<position>45.5,-23.5</position>
<gparam>LABEL_TEXT Q1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>85</ID>
<type>AA_LABEL</type>
<position>55.5,-23.5</position>
<gparam>LABEL_TEXT Q0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55.5,-40.5,55.5,-27</points>
<connection>
<GID>19</GID>
<name>N_in2</name></connection>
<intersection>-40.5 1</intersection>
<intersection>-33 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54,-40.5,55.5,-40.5</points>
<connection>
<GID>44</GID>
<name>OUT_0</name></connection>
<intersection>55.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>55.5,-33,65,-33</points>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<intersection>55.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>11,-49.5,48,-49.5</points>
<connection>
<GID>29</GID>
<name>OUT_0</name></connection>
<intersection>18.5 7</intersection>
<intersection>28 6</intersection>
<intersection>38.5 4</intersection>
<intersection>48 8</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>38.5,-49.5,38.5,-43.5</points>
<intersection>-49.5 1</intersection>
<intersection>-43.5 15</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>28,-49.5,28,-43.5</points>
<connection>
<GID>37</GID>
<name>clock</name></connection>
<intersection>-49.5 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>18.5,-49.5,18.5,-43.5</points>
<connection>
<GID>33</GID>
<name>clock</name></connection>
<intersection>-49.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>48,-49.5,48,-43.5</points>
<connection>
<GID>44</GID>
<name>clock</name></connection>
<intersection>-49.5 1</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>38.5,-43.5,40,-43.5</points>
<connection>
<GID>40</GID>
<name>clock</name></connection>
<intersection>38.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21.5,-56,21.5,-46.5</points>
<connection>
<GID>33</GID>
<name>clear</name></connection>
<intersection>-56 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>11.5,-56,51,-56</points>
<connection>
<GID>27</GID>
<name>OUT_0</name></connection>
<intersection>21.5 0</intersection>
<intersection>31 6</intersection>
<intersection>43 3</intersection>
<intersection>51 5</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>43,-56,43,-46.5</points>
<connection>
<GID>40</GID>
<name>clear</name></connection>
<intersection>-56 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>51,-56,51,-46.5</points>
<connection>
<GID>44</GID>
<name>clear</name></connection>
<intersection>-56 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>31,-56,31,-46.5</points>
<connection>
<GID>37</GID>
<name>clear</name></connection>
<intersection>-56 1</intersection></vsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46,-40.5,46,-27.5</points>
<connection>
<GID>40</GID>
<name>OUT_0</name></connection>
<connection>
<GID>15</GID>
<name>N_in2</name></connection>
<intersection>-40.5 5</intersection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>46,-32,65,-32</points>
<connection>
<GID>3</GID>
<name>IN_1</name></connection>
<intersection>46 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>46,-40.5,48,-40.5</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>46 0</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-40.5,35.5,-27</points>
<connection>
<GID>11</GID>
<name>N_in2</name></connection>
<intersection>-40.5 3</intersection>
<intersection>-40.5 3</intersection>
<intersection>-31 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>35.5,-31,65,-31</points>
<connection>
<GID>3</GID>
<name>IN_2</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>34,-40.5,40,-40.5</points>
<connection>
<GID>37</GID>
<name>OUT_0</name></connection>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-40.5,25,-27</points>
<connection>
<GID>7</GID>
<name>N_in2</name></connection>
<intersection>-40.5 1</intersection>
<intersection>-40.5 1</intersection>
<intersection>-30 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24.5,-40.5,28,-40.5</points>
<connection>
<GID>33</GID>
<name>OUT_0</name></connection>
<connection>
<GID>37</GID>
<name>IN_0</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25,-30,65,-30</points>
<connection>
<GID>3</GID>
<name>IN_3</name></connection>
<intersection>25 0</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>11.5,-40.5,18.5,-40.5</points>
<connection>
<GID>71</GID>
<name>OUT_0</name></connection>
<intersection>18.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>18.5,-40.5,18.5,-40.5</points>
<connection>
<GID>33</GID>
<name>IN_0</name></connection>
<intersection>-40.5 1</intersection></vsegment></shape></wire></page 1>
<page 2>
<PageViewport>-3.18452e-006,0,93.6,-90.8</PageViewport></page 2>
<page 3>
<PageViewport>-3.18452e-006,0,93.6,-90.8</PageViewport></page 3>
<page 4>
<PageViewport>-3.18452e-006,0,93.6,-90.8</PageViewport></page 4>
<page 5>
<PageViewport>-3.18452e-006,0,93.6,-90.8</PageViewport></page 5>
<page 6>
<PageViewport>-3.18452e-006,0,93.6,-90.8</PageViewport></page 6>
<page 7>
<PageViewport>-3.18452e-006,0,93.6,-90.8</PageViewport></page 7>
<page 8>
<PageViewport>-3.18452e-006,0,93.6,-90.8</PageViewport></page 8>
<page 9>
<PageViewport>-3.18452e-006,0,93.6,-90.8</PageViewport></page 9></circuit>